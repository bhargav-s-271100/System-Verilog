class transactor;
  randc bit [3:0]a,b;
  randc bit cin;
  bit valid;
  bit [4:0] c;
endclass
